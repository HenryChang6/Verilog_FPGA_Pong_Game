module state_machine(
    input  clk,
    input  rst,
    input  start,
    input  up1,
    input  up2,
    input  down1,
    input  down2,
    input  sec1, // ???
    output ball_x,
    output ball_y,
    output paddle1_x,
    output paddle1_y,
    output paddle2_x,
    output paddle2_y,
 );

 

endmodule