module test (clk, reset, red, green, blue, Hsync, Vsync, in, led, switch);
input clk, reset;
input switch;
output Hsync, Vsync;
output [3:0] led;
output [2:0] in;
output [3:0] red, green, blue;
wire [3:0] I_red, I_green, I_blue;
wire clk_div, active;
wire flag;
wire [11:0] v_cnt;
wire [11:0] h_cnt;
wire  [11:0] paddle;
wire [3:0] cnt;
FrequencyDivider u_FreqDiv(.clk(clk), .reset(reset), .clk_div(clk_div));
//RGBAdder u_Radder(.clk(clk_div), .reset(reset), .color(I_red), .button(switch));
//RGBAdder u_Gadder(.clk(clk_div), .reset(reset), .color(I_green), .button(switch));
RGBAdder adder(.clk(clk_div), .reset(reset), .color(cnt), .button(switch));
Graphic_gener(.paddle_1(paddle), .paddle_2(paddle), .ball_x(paddle), .ball_y(paddle), .v_cnt(v_cnt), .h_cnt(h_cnt), .flag(flag), .red(red), .green(green), .blue(blue));
vga_driver(.I_clk(clk), .I_rst_n(reset),.O_hs(Hsync),.O_vs(Vsync), .flag(flag), .v_cnt(v_cnt), .h_cnt(h_cnt));
assign led = cnt;
assign paddle[8:5] = cnt;
endmodule
