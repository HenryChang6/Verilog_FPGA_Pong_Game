module key_pad_controller (
    input clk, //100Hz
    input rst,
    input [3:0] kp_row,
    input [3:0] kp_col, 
    output up1, // A being pressed
    output up2, // 8 being pressed
    output down1, // 0 being pressed
    output down2, // 7 being pressed
);



endmodule