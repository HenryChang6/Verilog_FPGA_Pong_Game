score_counter sc(
    // input 
    .ball_x(ball_x),
    .ball_y(ball_y),
    // output
    .score1(score1),
    .score2(score2),
);

module score_counter(
    input ball_x,
    output score1,
    output score2,
);

endmodule